module converter_v (
    input  x2, x4, x8, x10, x20, z,
    output y2, y4, y8, y16, y32
);

    assign y2  = (z == 1'b0) ? 1'b1 : 
                 (~x20 & ~x10 & ~x8 & ~x4 & x2) |
                 (~x20 & ~x10 & ~x8 & x4 & x2) |
                 (~x20 & x10 & ~x8 & ~x4 & ~x2) |
                 (~x20 & x10 & ~x8 & x4 & ~x2) |
                 (~x20 & x10 & x8 & ~x4 & ~x2) |
                 (x20 & ~x10 & ~x8 & ~x4 & x2) |
                 (x20 & ~x10 & ~x8 & x4 & x2) |
                 (x20 & x10 & ~x8 & ~x4 & ~x2) |
                 (x20 & x10 & ~x8 & x4 & ~x2) |
                 (x20 & x10 & x8 & ~x4 & ~x2);

    assign y4  = (z == 1'b0) ? 1'b1 : 
                 (~x20 & ~x10 & ~x8 & x4 & ~x2) |
                 (~x20 & ~x10 & ~x8 & x4 & x2) |
                 (~x20 & x10 & ~x8 & ~x4 & x2) |
                 (~x20 & x10 & ~x8 & x4 & ~x2) |
                 (x20 & ~x10 & ~x8 & ~x4 & ~x2) |
                 (x20 & ~x10 & ~x8 & ~x4 & x2) |
                 (x20 & ~x10 & x8 & ~x4 & ~x2) |
                 (x20 & x10 & ~x8 & ~x4 & ~x2) |
                 (x20 & x10 & ~x8 & x4 & x2) |
                 (x20 & x10 & x8 & ~x4 & ~x2);

    assign y8  = (z== 1'b0) ? 1'b1 : 
                 (~x20 & ~x10 & x8 & ~x4 & ~x2) |
                 (~x20 & x10 & ~x8 & ~x4 & ~x2) |
                 (~x20 & x10 & ~x8 & ~x4 & x2) |
                 (~x20 & x10 & ~x8 & x4 & ~x2) |
                 (x20 & ~x10 & ~x8 & x4 & ~x2) |
                 (x20 & ~x10 & ~x8 & x4 & x2) |
                 (x20 & ~x10 & x8 & ~x4 & ~x2) |
                 (x20 & x10 & ~x8 & ~x4 & ~x2);

    assign y16 = (z== 1'b0) ? 1'b1 : 
                 (~x20 & x10 & ~x8 & x4 & x2) |
                 (~x20 & x10 & x8 & ~x4 & ~x2) |
                 (x20 & ~x10 & ~x8 & ~x4 & ~x2) |
                 (x20 & ~x10 & ~x8 & ~x4 & x2) |
                 (x20 & ~x10 & ~x8 & x4 & ~x2) |
                 (x20 & ~x10 & ~x8 & x4 & x2) |
                 (x20 & ~x10 & x8 & ~x4 & ~x2) |
                 (x20 & x10 & ~x8 & ~x4 & ~x2);

    assign y32 = (z== 1'b0) ? 1'b1 : 
                 (x20 & x10 & ~x8 & ~x4 & x2) |
                 (x20 & x10 & ~x8 & x4 & ~x2) |
                 (x20 & x10 & ~x8 & x4 & x2) |
                 (x20 & x10 & x8 & ~x4 & ~x2);

endmodule
